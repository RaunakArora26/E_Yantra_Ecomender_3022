
// instr_mem.v - instruction memory

module instr_mem #(parameter DATA_WIDTH = 32, ADDR_WIDTH = 32, MEM_SIZE = 512) (
    input       [ADDR_WIDTH-1:0] instr_addr,
    output      [DATA_WIDTH-1:0] instr
);

// array of 64 32-bit words or instructions
reg [DATA_WIDTH-1:0] instr_ram [0:MEM_SIZE-1];

// initial begin
//     // $readmemh("rv32i_test.hex", instr_ram);
// end
// Hardcoded Verilog Initialization
initial begin
  instr_ram[0] = 32'h02000117;
  instr_ram[1] = 32'h04010113;
  instr_ram[2] = 32'h02000197;
  instr_ram[3] = 32'h7F818193;
  instr_ram[4] = 32'h02000517;
  instr_ram[5] = 32'hFF050513;
  instr_ram[6] = 32'h33800593;
  instr_ram[7] = 32'h00000613;
  instr_ram[8] = 32'h2D8000EF;
  instr_ram[9] = 32'h02000517;
  instr_ram[10] = 32'hFDC50513;
  instr_ram[11] = 32'h00000593;
  instr_ram[12] = 32'h00000613;
  instr_ram[13] = 32'h2E8000EF;
  instr_ram[14] = 32'h02000517;
  instr_ram[15] = 32'hFC850513;
  instr_ram[16] = 32'h2B0000EF;
  instr_ram[17] = 32'h00000513;
  instr_ram[18] = 32'h00000593;
  instr_ram[19] = 32'h008000EF;
  instr_ram[20] = 32'h0000006F;
  instr_ram[21] = 32'hFF010113;
  instr_ram[22] = 32'h00112623;
  instr_ram[23] = 32'h00812423;
  instr_ram[24] = 32'h00001737;
  instr_ram[25] = 32'h02000437;
  instr_ram[26] = 32'h44200793;
  instr_ram[27] = 32'h00F42823;
  instr_ram[28] = 32'h80570793;
  instr_ram[29] = 32'h00F42A23;
  instr_ram[30] = 32'h03A00793;
  instr_ram[31] = 32'h00F42C23;
  instr_ram[32] = 32'h00400793;
  instr_ram[33] = 32'h00F42E23;
  instr_ram[34] = 32'h02F42023;
  instr_ram[35] = 32'h02F42223;
  instr_ram[36] = 32'h38100793;
  instr_ram[37] = 32'h02F42423;
  instr_ram[38] = 32'h04000793;
  instr_ram[39] = 32'h02F42623;
  instr_ram[40] = 32'h02F42823;
  instr_ram[41] = 32'h02F42A23;
  instr_ram[42] = 32'h050017B7;
  instr_ram[43] = 32'h80178793;
  instr_ram[44] = 32'h02F42C23;
  instr_ram[45] = 32'h000817B7;
  instr_ram[46] = 32'h40278793;
  instr_ram[47] = 32'h02F42E23;
  instr_ram[48] = 32'h000077B7;
  instr_ram[49] = 32'h80078793;
  instr_ram[50] = 32'h04F42023;
  instr_ram[51] = 32'h000197B7;
  instr_ram[52] = 32'h04F42423;
  instr_ram[53] = 32'h000047B7;
  instr_ram[54] = 32'h04F42623;
  instr_ram[55] = 32'h000647B7;
  instr_ram[56] = 32'h04F42823;
  instr_ram[57] = 32'h000107B7;
  instr_ram[58] = 32'h04F42A23;
  instr_ram[59] = 32'h002907B7;
  instr_ram[60] = 32'h04F42C23;
  instr_ram[61] = 32'h001417B7;
  instr_ram[62] = 32'h80078793;
  instr_ram[63] = 32'h04F42E23;
  instr_ram[64] = 32'h000807B7;
  instr_ram[65] = 32'h06F42023;
  instr_ram[66] = 32'h00C407B7;
  instr_ram[67] = 32'h06F42223;
  instr_ram[68] = 32'h002007B7;
  instr_ram[69] = 32'h06F42423;
  instr_ram[70] = 32'h412007B7;
  instr_ram[71] = 32'h06F42623;
  instr_ram[72] = 32'h028007B7;
  instr_ram[73] = 32'h40078793;
  instr_ram[74] = 32'h06F42823;
  instr_ram[75] = 32'h010007B7;
  instr_ram[76] = 32'h06F42A23;
  instr_ram[77] = 32'h180007B7;
  instr_ram[78] = 32'h40078793;
  instr_ram[79] = 32'h06F42C23;
  instr_ram[80] = 32'h040007B7;
  instr_ram[81] = 32'h06F42E23;
  instr_ram[82] = 32'h640007B7;
  instr_ram[83] = 32'h08F42023;
  instr_ram[84] = 32'h100007B7;
  instr_ram[85] = 32'h04E42223;
  instr_ram[86] = 32'h08F42223;
  instr_ram[87] = 32'h908007B7;
  instr_ram[88] = 32'h08F42423;
  instr_ram[89] = 32'h400007B7;
  instr_ram[90] = 32'h08F42623;
  instr_ram[91] = 32'h02000613;
  instr_ram[92] = 32'h02800593;
  instr_ram[93] = 32'h0D040513;
  instr_ram[94] = 32'h1A4000EF;
  instr_ram[95] = 32'h0FF00593;
  instr_ram[96] = 32'h0B140513;
  instr_ram[97] = 32'h02000613;
  instr_ram[98] = 32'h194000EF;
  instr_ram[99] = 32'h00044783;
  instr_ram[100] = 32'h020005B7;
  instr_ram[101] = 32'hFA000537;
  instr_ram[102] = 32'h0FF7F793;
  instr_ram[103] = 32'h00F40433;
  instr_ram[104] = 32'h0C040823;
  instr_ram[105] = 32'h01F00793;
  instr_ram[106] = 32'hCD050513;
  instr_ram[107] = 32'h00100E13;
  instr_ram[108] = 32'h02800F93;
  instr_ram[109] = 32'h0D058293;
  instr_ram[110] = 32'h02000E93;
  instr_ram[111] = 32'h0F058F13;
  instr_ram[112] = 32'h0D058713;
  instr_ram[113] = 32'h0480006F;
  instr_ram[114] = 32'h00082303;
  instr_ram[115] = 32'h00DE1633;
  instr_ram[116] = 32'h00667633;
  instr_ram[117] = 32'h02060463;
  instr_ram[118] = 32'h00074603;
  instr_ram[119] = 32'h03F60063;
  instr_ram[120] = 32'h00568333;
  instr_ram[121] = 32'h00034383;
  instr_ram[122] = 32'h00160613;
  instr_ram[123] = 32'h00765863;
  instr_ram[124] = 32'h00C30023;
  instr_ram[125] = 32'h00D58633;
  instr_ram[126] = 32'h0B1608A3;
  instr_ram[127] = 32'h00168693;
  instr_ram[128] = 32'hFDD694E3;
  instr_ram[129] = 32'h00170713;
  instr_ram[130] = 32'h01E70E63;
  instr_ram[131] = 32'h03070893;
  instr_ram[132] = 32'h00271813;
  instr_ram[133] = 32'h0FF8F893;
  instr_ram[134] = 32'h00A80833;
  instr_ram[135] = 32'h00000693;
  instr_ram[136] = 32'hFA9FF06F;
  instr_ram[137] = 32'hFFF78793;
  instr_ram[138] = 32'h0FF7F793;
  instr_ram[139] = 32'hF8079AE3;
  instr_ram[140] = 32'h02000737;
  instr_ram[141] = 32'h00474703;
  instr_ram[142] = 32'h020006B7;
  instr_ram[143] = 32'h00000613;
  instr_ram[144] = 32'h0FF77713;
  instr_ram[145] = 32'h0FF00593;
  instr_ram[146] = 32'h0B168513;
  instr_ram[147] = 32'h04B71663;
  instr_ram[148] = 32'hFFF60693;
  instr_ram[149] = 32'h02000737;
  instr_ram[150] = 32'h0FF6F693;
  instr_ram[151] = 32'h0EF70713;
  instr_ram[152] = 32'h04D7EA63;
  instr_ram[153] = 32'h00070793;
  instr_ram[154] = 32'h020006B7;
  instr_ram[155] = 32'h01178713;
  instr_ram[156] = 32'h0FF77713;
  instr_ram[157] = 32'h06C76663;
  instr_ram[158] = 32'h020007B7;
  instr_ram[159] = 32'h00100713;
  instr_ram[160] = 32'h00E78623;
  instr_ram[161] = 32'h00C12083;
  instr_ram[162] = 32'h00812403;
  instr_ram[163] = 32'h00000513;
  instr_ram[164] = 32'h01010113;
  instr_ram[165] = 32'h00008067;
  instr_ram[166] = 32'h00160813;
  instr_ram[167] = 32'h00C68633;
  instr_ram[168] = 32'h0EE607A3;
  instr_ram[169] = 32'h00A70733;
  instr_ram[170] = 32'h00074703;
  instr_ram[171] = 32'h0FF87613;
  instr_ram[172] = 32'hF9DFF06F;
  instr_ram[173] = 32'h00E685B3;
  instr_ram[174] = 32'h00E78533;
  instr_ram[175] = 32'h0005C883;
  instr_ram[176] = 32'h00054803;
  instr_ram[177] = 32'h00178793;
  instr_ram[178] = 32'h01150023;
  instr_ram[179] = 32'hFFF68693;
  instr_ram[180] = 32'h01058023;
  instr_ram[181] = 32'h0FF7F793;
  instr_ram[182] = 32'h0FF6F693;
  instr_ram[183] = 32'hF85FF06F;
  instr_ram[184] = 32'h0007C703;
  instr_ram[185] = 32'h00178793;
  instr_ram[186] = 32'h00E68423;
  instr_ram[187] = 32'hF81FF06F;
  instr_ram[188] = 32'h00050213;
  instr_ram[189] = 32'h00008067;
  instr_ram[190] = 32'h00050313;
  instr_ram[191] = 32'h00060E63;
  instr_ram[192] = 32'h00058383;
  instr_ram[193] = 32'h00730023;
  instr_ram[194] = 32'hFFF60613;
  instr_ram[195] = 32'h00130313;
  instr_ram[196] = 32'h00158593;
  instr_ram[197] = 32'hFE0616E3;
  instr_ram[198] = 32'h00008067;
  instr_ram[199] = 32'h00050313;
  instr_ram[200] = 32'h00060A63;
  instr_ram[201] = 32'h00B30023;
  instr_ram[202] = 32'hFFF60613;
  instr_ram[203] = 32'h00130313;
  instr_ram[204] = 32'hFE061AE3;
  instr_ram[205] = 32'h00008067;
  instr_ram[206] = 32'h00000000;
  instr_ram[207] = 32'h00000000;
  instr_ram[208] = 32'h00000000;
  instr_ram[209] = 32'h00000000;
  instr_ram[210] = 32'h00000000;
  instr_ram[211] = 32'h00000000;
  instr_ram[212] = 32'h00000000;
  instr_ram[213] = 32'h00000000;
  instr_ram[214] = 32'h00000000;
  instr_ram[215] = 32'h00000000;
  instr_ram[216] = 32'h00000000;
  instr_ram[217] = 32'h00000000;
  instr_ram[218] = 32'h00000000;
  instr_ram[219] = 32'h00000000;
  instr_ram[220] = 32'h00000000;
  instr_ram[221] = 32'h00000000;
  instr_ram[222] = 32'h00000000;
  instr_ram[223] = 32'h00000000;
  instr_ram[224] = 32'h00000000;
  instr_ram[225] = 32'h00000000;
  instr_ram[226] = 32'h00000000;
  instr_ram[227] = 32'h00000000;
  instr_ram[228] = 32'h00000000;
  instr_ram[229] = 32'h00000000;
  instr_ram[230] = 32'h00000000;
  instr_ram[231] = 32'h00000000;
  instr_ram[232] = 32'h00000000;
  instr_ram[233] = 32'h00000000;
  instr_ram[234] = 32'h00000000;
  instr_ram[235] = 32'h00000000;
  instr_ram[236] = 32'h00000000;
  instr_ram[237] = 32'h00000000;
  instr_ram[238] = 32'h00000000;
  instr_ram[239] = 32'h00000000;
  instr_ram[240] = 32'h00000000;
  instr_ram[241] = 32'h00000000;
  instr_ram[242] = 32'h00000000;
  instr_ram[243] = 32'h00000000;
  instr_ram[244] = 32'h00000000;
  instr_ram[245] = 32'h00000000;
  instr_ram[246] = 32'h00000000;
  instr_ram[247] = 32'h00000000;
  instr_ram[248] = 32'h00000000;
  instr_ram[249] = 32'h00000000;
  instr_ram[250] = 32'h00000000;
  instr_ram[251] = 32'h00000000;
  instr_ram[252] = 32'h00000000;
  instr_ram[253] = 32'h00000000;
  instr_ram[254] = 32'h00000000;
  instr_ram[255] = 32'h00000000;
end


// word-aligned memory access
// combinational read logic
assign instr = instr_ram[instr_addr[31:2]];

endmodule

